`include "CPU_Defines.v"

`timescale 1ns/1ns

module CPU_Registers (
	input i_reset,
	input i_clock,

	input i_read,
	input [4:0] i_read_rs1_idx,
	input [4:0] i_read_rs2_idx,
	output [31:0] o_rs1,
	output [31:0] o_rs2,

	input i_write,
	input [4:0] i_write_rd_idx,
	input [31:0] i_rd
);
	assign o_rs1 = rs1;
	assign o_rs2 = rs2;

	reg [31:0] r[31:0];
	reg [31:0] rs1 = 0;
	reg [31:0] rs2 = 0;

    initial begin
        r[ 0] = 32'h0000_0000;
        r[ 1] = 32'h0000_0000;
        r[ 2] = 32'h1000_0400 - 4;	// sp	
        r[ 3] = 32'h0000_0000;
        r[ 4] = 32'h0000_0000;
        r[ 5] = 32'h0000_0000;
        r[ 6] = 32'h0000_0000;
        r[ 7] = 32'h0000_0000;
        r[ 8] = 32'h0000_0000;
        r[ 9] = 32'h0000_0000;
        r[10] = 32'h0000_0000;
        r[11] = 32'h0000_0000;
        r[12] = 32'h0000_0000;
        r[13] = 32'h0000_0000;
        r[14] = 32'h0000_0000;
        r[15] = 32'h0000_0000;
        r[16] = 32'h0000_0000;
        r[17] = 32'h0000_0000;
        r[18] = 32'h0000_0000;
        r[19] = 32'h0000_0000;
        r[20] = 32'h0000_0000;
        r[21] = 32'h0000_0000;
        r[22] = 32'h0000_0000;
        r[23] = 32'h0000_0000;
        r[24] = 32'h0000_0000;
        r[25] = 32'h0000_0000;
        r[26] = 32'h0000_0000;
        r[27] = 32'h0000_0000;
        r[28] = 32'h0000_0000;
        r[29] = 32'h0000_0000;
        r[30] = 32'h0000_0000;
        r[31] = 32'h0000_0000;       
    end

	always @(posedge i_clock, posedge i_reset)
	begin
		if (i_reset) begin
			rs1 <= 0;
			rs2 <= 0;

			r[ 0] <= 32'h0000_0000;
			r[ 1] <= 32'h0000_0000;
			r[ 2] <= 32'h1000_0400 - 4;	// sp	
			r[ 3] <= 32'h0000_0000;
			r[ 4] <= 32'h0000_0000;
			r[ 5] <= 32'h0000_0000;
			r[ 6] <= 32'h0000_0000;
			r[ 7] <= 32'h0000_0000;
			r[ 8] <= 32'h0000_0000;
			r[ 9] <= 32'h0000_0000;
			r[10] <= 32'h0000_0000;
			r[11] <= 32'h0000_0000;
			r[12] <= 32'h0000_0000;
			r[13] <= 32'h0000_0000;
			r[14] <= 32'h0000_0000;
			r[15] <= 32'h0000_0000;
			r[16] <= 32'h0000_0000;
			r[17] <= 32'h0000_0000;
			r[18] <= 32'h0000_0000;
			r[19] <= 32'h0000_0000;
			r[20] <= 32'h0000_0000;
			r[21] <= 32'h0000_0000;
			r[22] <= 32'h0000_0000;
			r[23] <= 32'h0000_0000;
			r[24] <= 32'h0000_0000;
			r[25] <= 32'h0000_0000;
			r[26] <= 32'h0000_0000;
			r[27] <= 32'h0000_0000;
			r[28] <= 32'h0000_0000;
			r[29] <= 32'h0000_0000;
			r[30] <= 32'h0000_0000;
			r[31] <= 32'h0000_0000;
		end
		else begin
			if (i_read) begin
                rs1 <= (i_read_rs1_idx != 0) ? r[i_read_rs1_idx] : 32'h0;
                rs2 <= (i_read_rs2_idx != 0) ? r[i_read_rs2_idx] : 32'h0;
			end
			if (i_write) begin
				r[i_write_rd_idx] <= i_rd;
			end
		end
	end

endmodule