
`timescale 1ns/1ns

module Timer (
	input i_reset,
	input i_clock,
	input i_request,
	input i_rw,
	input [3:0] i_address,
	input [31:0] i_wdata,
	output bit [31:0] o_rdata,
	output bit o_ready,

	output bit o_interrupt
);

	bit [63:0] cycles = 0;
	bit [63:0] compare = { 64{1'b1} };
	bit request = 0;

	initial begin
		o_ready = 1'b0;
		o_interrupt = 1'b0;
	end

	always_ff @(posedge i_clock) begin
		if (i_reset) begin
			cycles <= 0;
		end
		else begin
			cycles <= cycles + 64'h1;
			o_interrupt <= ((cycles == compare) ? 1'b1 : 1'b0);
		end
	end

	always_ff @(posedge i_clock) begin
		request <= i_request;
		if (i_request && !request) begin
			if (!i_rw) begin
				case (i_address)
					4'h0: o_rdata <= cycles[31:0];
					4'h1: o_rdata <= cycles[63:32];
					4'h2: o_rdata <= compare[31:0];
					4'h3: o_rdata <= compare[63:32];
					default: o_rdata <= 0;
				endcase
			end
			else begin
				case (i_address)
					4'h2: compare[31:0] <= i_wdata;
					4'h3: compare[63:32] <= i_wdata;
					default:;
				endcase
			end
			o_ready <= 1;
		end
		else if (!i_request)
			o_ready <= 0;
	end
	
endmodule
