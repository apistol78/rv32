`include "CPU_Defines.sv"

`timescale 1ns/1ns

module CPU_Decode(
	input wire i_reset,
	input wire i_clock,
	output reg o_fault,

	// Input
	output o_busy,
	input fetch_data_t i_data,
	
	// Output
	input i_execute_busy,
	output decode_data_t o_data
);

	`include "Instructions_ops.sv"

	`undef INSTRUCTION
	`define INSTRUCTION i_data.instruction
	`include "Instructions_decode.sv"
	
	// Alias symbols for generated code.
	`undef ZERO
	`undef RS1
	`undef RS2
	`undef PC
	`undef IMM
	`define ZERO 3'd0
	`define RS1 3'd1
	`define RS2 3'd2
	`define PC	3'd3
	`define IMM 3'd4
	`include "Instructions_alu.sv"

	`include "Instructions_memory.sv"

	wire [31:0] inst_B_imm = { { 20{ `INSTRUCTION[31] } }, `INSTRUCTION[7], `INSTRUCTION[30:25], `INSTRUCTION[11:8], 1'b0 };
	wire [31:0] inst_I_imm = { { 21{ `INSTRUCTION[31] } }, `INSTRUCTION[30:20] };
	wire [31:0] inst_J_imm = { { 12{ `INSTRUCTION[31] } }, `INSTRUCTION[19:12], `INSTRUCTION[20], `INSTRUCTION[30:21], 1'b0 };
	wire [31:0] inst_S_imm = { { 21{ `INSTRUCTION[31] } }, `INSTRUCTION[30:25], `INSTRUCTION[11:7] };
	wire [31:0] inst_U_imm = { `INSTRUCTION[31:12], 12'b0 };
	wire [31:0] inst_R_imm = { 26'b0, `INSTRUCTION[25:20] };
	wire [31:0] inst_CSR_imm = { 20'b0, `INSTRUCTION[31:20] };
	
	wire have_RS1 = is_B | is_I | is_R | is_S | is_CSR;
	wire have_RS2 = is_B | is_R | is_S;
	wire have_RD  = is_I | is_J | is_R | is_U | is_CSR;

	decode_data_t dataC = 0;
	decode_data_t dataN = 0;

	assign o_busy = i_execute_busy;
	assign o_data = !i_execute_busy ? dataC : dataN;

	initial begin
		o_fault = 0;
	end

	always_ff @(posedge i_clock) begin
		if (!i_execute_busy)
			dataN <= dataC;
	end

	always_ff @(posedge i_clock) begin
		if (i_reset) begin
			dataC <= 0;
			dataN <= 0;
			o_fault <= 0;
		end
		else begin

			if (i_data.tag != dataC.tag) begin

				dataC.instruction <= i_data.instruction;
				dataC.pc <= i_data.pc;

				dataC.inst_rs1 <= have_RS1 ? `INSTRUCTION[19:15] : 5'h0;
				dataC.inst_rs2 <= have_RS2 ? `INSTRUCTION[24:20] : 5'h0;
				dataC.inst_rd  <= have_RD  ? `INSTRUCTION[ 11:7] : 5'h0;
				
				dataC.imm <=
					is_B ? inst_B_imm :
					is_I ? inst_I_imm :
					is_J ? inst_J_imm :
					is_S ? inst_S_imm :
					is_U ? inst_U_imm :
					is_R ? inst_R_imm :
					is_CSR ? inst_CSR_imm :
					32'h0;
				
				dataC.arithmetic <= is_ARITHMETIC;
				dataC.compare <= is_COMPARE;
				dataC.complx <= is_COMPLEX;
				dataC.jump <= is_JUMP;
				dataC.jump_conditional <= is_JUMP_CONDITIONAL;

				dataC.alu_operation <= alu_operation;
				dataC.alu_operand1 <= alu_operand1;
				dataC.alu_operand2 <= alu_operand2;

				dataC.memory_read <= memory_read;
				dataC.memory_write <= memory_write;
				dataC.memory_width <= memory_width;
				dataC.memory_signed <= memory_signed;
				
				`define OP dataC.op
				`include "Instructions_decode_ops.sv"

				if (is_ARITHMETIC || is_COMPARE || is_COMPLEX || is_JUMP || is_JUMP_CONDITIONAL || is_MEMORY) begin
					dataC.tag <= i_data.tag;
				end
				else begin
					// Invalid or unsupported instructions end here.
					o_fault <= 1;
				end
			end
		end
	end

endmodule
